<?php

	/*****************************************************************************

		The Swedish nls files are contributed by: Niklas Koskela <ntkk@htc.se>
                                                      Karl Thysell <karl@htc.se>

	*****************************************************************************/

	$ARnls["xp_new"]						=	"L&auml;gg till nytt objekt";
	$ARnls["xp_rename"]						=	"Byt namn ";
	$ARnls["xp_copy"]						=	"Kopiera ";
	$ARnls["xp_link"]						=	"L&auml;nk ";
	$ARnls["xp_edit"]						=	"&auml;ndra ";
	$ARnls["xp_shortcut"]					=	"&auml;ndra genv&auml;g";
	$ARnls["xp_delete"]						=	"Radera ";
	$ARnls["xp_cache"]						=	"S&auml;tt cache f&ouml;r ";
	$ARnls["xp_templates"]					=	"S&auml;tt mallar f&ouml;r ";
	$ARnls["xp_customfields"]				=	"S&auml;tt anpassade f&auml;lt f&ouml;r ";
	$ARnls["xp_language"]					=	"S&auml;tt spr&aring;k f&ouml;r ";
	$ARnls["xp_grants"]						=	"S&auml;tt r&auml;ttigheter f&ouml;r ";
	$ARnls["xp_types"]						=	"S&auml;tt typtr&auml;d f&ouml;r ";
	$ARnls["xp_priority"]					=	"S&auml;tt prioritet f&ouml;r ";
	$ARnls["xp_viewweb"]					=	"Visa webbsida ";
	$ARnls["xp_view"]						=	"Visa";
	$ARnls["xp_explore"]					=	"Utforska";
	
	//headers
	$ARnls["xp_settings"]					=	"Inst&auml;llningar";
	$ARnls["xp_info"]						=	"Information";
	$ARnls["xp_detailsH"]					=	"Mera...";
	$ARnls["xp_browsebyletter"]				=	"Bl&auml;ddra per bokstav";
	$ARnls["xp_browsebydate"]				=	"Bl&auml;ddra per datum";
	
	//toolbar
	$ARnls["xp_up"]							= 	"Upp";
	$ARnls["xp_search"]						= 	"S&ouml;k";
	$ARnls["xp_folders"]					= 	"Mappar";
	$ARnls["xp_small"]						= 	"Lista";
	$ARnls["xp_large"]						= 	"Ikoner";
	$ARnls["xp_details"]					= 	"Detaljer";
	$ARnls["xp_iconview"]					= 	"V&auml;lj Ikon-vy";
	$ARnls["xp_import"]						= 	"Importera";
	$ARnls["xp_export"]						= 	"Exportera";
	$ARnls["xp_preferences"]				= 	"Egenskaper";
	$ARnls["xp_help"]						= 	"Hj&auml;lp";
	$ARnls["xp_tutorials"]					= 	"V&auml;gledning";
	$ARnls["xp_about"]						= 	"Om...";


?>
