<?php

	/*****************************************************************************

		The Swedish nls files are contributed by: Niklas Koskela <ntkk@htc.se>
                                                      Karl Thysell <karl@htc.se>

	*****************************************************************************/

	// Attention: The WYSIWYG editor and its context menus require UTF-8!
	// (The external dialogs do not)

	// lib/widgets/htmledit/ie/edit.php

	$ARnls["e_cut"]				=	"Klipp ut";
	$ARnls["e_copy"]			=	"Kopiera";
	$ARnls["e_paste"]			=	"Klistra in";
	$ARnls["e_delete"]			=	"Radera";

	$ARnls["e_insertrow"]			=	"Infoga Rader";
	$ARnls["e_deleterows"]			=	"Radera Rader";
	$ARnls["e_insertcol"]			=	"Infoga Kolumner";
	$ARnls["e_deletecols"]			=	"Raders Kolumner";
	$ARnls["e_insertcell"]			=	"Infoga Celler";
	$ARnls["e_deletecells"]			=	"Raders Celler";
	$ARnls["e_mergecells"]			=	"Sammanfoga Celler";
	$ARnls["e_splitcell"]			=	"Dela Celler";

	$ARnls["e_z_order"]			=	"Z Order";
	$ARnls["e_send_to_back"]		=	"S&auml;nd L&auml;ngst Bak";
	$ARnls["e_bring_to_front"]		=	"S&auml;nd L&auml;ngst Fram";
	$ARnls["e_send_backward"]		=	"S&auml;nd Bak&aring;t";
	$ARnls["e_bring_forward"]		=	"S&auml;nd Fram&aring;t";
	$ARnls["e_send_below_text"]		=	"S&auml;nd Under Text";
	$ARnls["e_bring_above_text"]		=	"S&auml;nd &ouml;ver Text";
	$ARnls["e_visible_borders"]		=	"Synliga Kanter";
	$ARnls["e_show_details"]		=	"Visa Detaljer";
	$ARnls["e_make_absolute"]		=	"G&ouml;r Absolut";
	$ARnls["e_lock"]			=	"L&aring;s";
	$ARnls["e_snap_to_grid"]		=	"F&auml;st Mot M&ouml;nster";

	$ARnls["e_file"]			=	"Fil";
	$ARnls["e_save_file"]			=	"Spara Fil";

	$ARnls["e_edit"]			=	"&Auml;ndra";
	$ARnls["e_undo"]			=	"&Aring;ngra";
	$ARnls["e_redo"]			=	"Upprepa";
	$ARnls["e_select_all"]			=	"Markera Allt";
	$ARnls["e_find"]			=	"S&ouml;k...";

	$ARnls["e_view"]			=	"Vy";
	$ARnls["e_standard"]			=	"Standard";
	$ARnls["e_toolbars"]			=	"Verktygsf&auml;lt";
	$ARnls["e_formatting"]			=	"Formatering";
	$ARnls["e_absolute_positioning"]	=	"Absolut Positionering";
	$ARnls["e_table"]			=	"Tabell";

	$ARnls["e_bold"]			=	"Fet";
	$ARnls["e_italic"]			=	"Kursiv";
	$ARnls["e_underline"]			=	"Understruken";

	$ARnls["e_set_foreground_color"]	=	"S&auml;tt F&ouml;rgrunds F&auml;rg...";
	$ARnls["e_set_background_color"]	=	"S&auml;tt Bakgrunds F&auml;rg...";
	$ARnls["e_foreground_color"]		=	"F&ouml;rgrunds F&auml;rg";
	$ARnls["e_background_color"]		=	"Bakgrunds F&auml;rg";

	$ARnls["e_align_left"]			=	"Justera V&auml;nster";
	$ARnls["e_align_center"]		=	"Centrera";
	$ARnls["e_align_right"]			=	"Justera H&ouml;ger";

	$ARnls["e_numbered_list"]		=	"Numrerad Lista";
	$ARnls["e_bulleted_list"]		=	"Punkt Lista";

	$ARnls["e_decrease_indent"]		=	"Minska Indrag";
	$ARnls["e_increase_indent"]		=	"&Ouml;ka Indrag";

	$ARnls["e_link"]			=	"L&auml;nk";
	$ARnls["e_insert_image"]		=	"Infoga Bild";
	$ARnls["e_insert_table"]		=	"Infoga Tabell";

	// lib/templates/pobject/edit.object.html.selectcolor.phtml

	$ARnls["e_select_color"]		=	"V&auml;lj F&auml;rg";
	$ARnls["e_color"]			=	"F&auml;rg";

	// lib/templates/pobject/edit.object.html.image.phtml

	$ARnls["e_picture"]			=	"Bild";
	$ARnls["e_picture_source"]		=	"Bild&nbsp;K&auml;lla";
	$ARnls["e_alternate_text"]		=	"Alternativ&nbsp;Text";
	$ARnls["e_layout"]			=	"Layout";
	$ARnls["e_alignment"]			=	"Placering";
	$ARnls["e_border_thickness"]		=	"Kant&nbsp;Tjocklek";
	$ARnls["e_spacing"]			=	"Mellanrum";
	$ARnls["e_horizontal"]			=	"Horisontell";
	$ARnls["e_vertical"]			=	"Vertikal";

	// lib/templates/pobject/edit.object.html.link*.phtml

	$ARnls["e_hyperlink"]			=	"Hyperl&auml;nk";
	$ARnls["e_hyperlink_information"]	=	"Hyperl&auml;nks&nbsp;Information";
	$ARnls["e_hyperlink_type"]		=	"Typ";
	$ARnls["e_hyperlink_path"]		=	"S&ouml;kv&auml;g";
	$ARnls["e_hyperlink_affiliate"]		=	"Anslut";

?>