<?PHP

	/*****************************************************************************

		The Swedish nls files are contributed by: Niklas Koskela <ntkk@htc.se>
                                                      Karl Thysell <karl@htc.se>

	*****************************************************************************/

	$ARnls["m_about"]						=	"Om&nbsp;Ariadne";
	$ARnls["m_cache"]						=	"Cache";
	$ARnls["m_config"]						=	"Konfiguration";
	$ARnls["m_copy"]						=	"Kopiera";
	$ARnls["m_custom"]						=	"Anpassade&nbsp;F&auml;lt";
	$ARnls["m_data"]						=	"Data";
	$ARnls["m_delete"]						=	"Ta bort";
	$ARnls["m_details"]						=	"Detaljer";
	$ARnls["m_edit"]						=	"Redigera";
	$ARnls["m_explorerbar"]					=	"Explorer&nbsp;F&auml;lt";
	$ARnls["m_export"]						=	"Exportera";
	$ARnls["m_find"]						=	"S&ouml;k";
	$ARnls["m_fonts"]						=	"Teckensnitt";
	$ARnls["m_grants"]						=	"R&auml;ttigheter";
	$ARnls["m_help"]						=	"Hj&auml;lp";
	$ARnls["m_import"]						=	"Importera";
	$ARnls["m_index"]						=	"Index";
	$ARnls["m_language"]					=	"Spr&aring;k";
	$ARnls["m_large"]						=	"Stora&nbsp;Ikoner";
	$ARnls["m_layout"]						=	"Layout";
	$ARnls["m_link"]						=	"L&auml;nk";
	$ARnls["m_logoff"]						=	"Logga&nbsp;av";
	$ARnls["m_new"]							=	"Nytt";
	$ARnls["m_object"]						=	"Objekt";
	$ARnls["m_preferences"]					=	"Inst&auml;llningar";
	$ARnls["m_priority"]					=	"Prioritet";
	$ARnls["m_rename"]						=	"Byt namn";
	$ARnls["m_search"]						=	"S&ouml;k";
	$ARnls["m_shortcut"]					=	"Genv&auml;g";
	$ARnls["m_small"]						=	"Sm&aring;&nbsp;Ikoner";
	$ARnls["m_templates"]					=	"Mallar";
	$ARnls["m_tutorials"]					=	"V&auml;gledning";
	$ARnls["m_types"]						=	"Typer";
	$ARnls["m_view"]						=	"Visa";
	$ARnls["m_web"]							=	"Webbsida";
	$ARnls["m_page"]						=	"Sida";
?>