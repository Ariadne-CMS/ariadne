<?php

	/*****************************************************************************

		The Swedish nls files are contributed by: Niklas Koskela <ntkk@htc.se>
                                                      Karl Thysell <karl@htc.se>

	*****************************************************************************/
	$ARnls["ariadne:about"]                         =    "Om...";
	$ARnls["ariadne:ace_editor"]                    =    "Ace Editor";
//	$ARnls["ariadne:apkg:depends_on"]               =    "Depends on"; // value from english
//	$ARnls["ariadne:apkg:install"]                  =    "Install"; // value from english
//	$ARnls["ariadne:apkg:install_package"]          =    "Install Ariadne package"; // value from english
//	$ARnls["ariadne:apkg:installing"]               =    "Installing Ariadne package..."; // value from english
//	$ARnls["ariadne:apkg:maintainer"]               =    "Maintainer"; // value from english
//	$ARnls["ariadne:apkg:package_information"]      =    "Package information"; // value from english
//	$ARnls["ariadne:apkg:target_location"]          =    "Package install location"; // value from english
//	$ARnls["ariadne:apkg:version"]                  =    "Version"; // value from english
//	$ARnls["ariadne:browse:select"]                 =    "Select"; // value from english
	$ARnls["ariadne:browsebydate"]                  =    "Bl&auml;ddra per datum";
	$ARnls["ariadne:browsebyletter"]                =    "Bl&auml;ddra per bokstav";
//	$ARnls["ariadne:browsetotarget"]                =    "Browse to target"; // value from english
//	$ARnls["ariadne:by"]                            =    "By"; // value from english
	$ARnls["ariadne:cache"]                         =    "S&auml;tt cache f&ouml;r ";
//	$ARnls["ariadne:change_priority"]               =    "Change priority"; // value from english
//	$ARnls["ariadne:childrenonly"]                  =    "Children only"; // value from english
//	$ARnls["ariadne:close"]                         =    "Close"; // value from english
	$ARnls["ariadne:copy"]                          =    "Kopiera ";
//	$ARnls["ariadne:created"]                       =    "Created"; // value from english
//	$ARnls["ariadne:currentandchildren"]            =    "Current object and children"; // value from english
//	$ARnls["ariadne:currentobjectonly"]             =    "Current object only"; // value from english
//	$ARnls["ariadne:currentowner"]                  =    "Current owner"; // value from english
	$ARnls["ariadne:customfields"]                  =    "S&auml;tt anpassade f&auml;lt f&ouml;r ";
	$ARnls["ariadne:delete"]                        =    "Radera ";
	$ARnls["ariadne:details"]                       =    "Detaljer";
	$ARnls["ariadne:detailsH"]                      =    "Mera...";
	$ARnls["ariadne:edit"]                          =    "&auml;ndra ";
//	$ARnls["ariadne:editor:align_absbottom"]        =    "Absbottom"; // value from english
//	$ARnls["ariadne:editor:align_absmiddle"]        =    "Absmiddle"; // value from english
//	$ARnls["ariadne:editor:align_baseline"]         =    "Baseline"; // value from english
//	$ARnls["ariadne:editor:align_bottom"]           =    "Bottom"; // value from english
//	$ARnls["ariadne:editor:align_left"]             =    "Left"; // value from english
//	$ARnls["ariadne:editor:align_middle"]           =    "Middle"; // value from english
//	$ARnls["ariadne:editor:align_not_set"]          =    "None"; // value from english
//	$ARnls["ariadne:editor:align_right"]            =    "Right"; // value from english
//	$ARnls["ariadne:editor:align_texttop"]          =    "Text top"; // value from english
//	$ARnls["ariadne:editor:align_top"]              =    "Top"; // value from english
//	$ARnls["ariadne:editor:alignment"]              =    "Alignment"; // value from english
//	$ARnls["ariadne:editor:anchor"]                 =    "Anchor"; // value from english
//	$ARnls["ariadne:editor:behaviour"]              =    "Behaviour"; // value from english
//	$ARnls["ariadne:editor:currentwindow"]          =    "Open in current window"; // value from english
//	$ARnls["ariadne:editor:external_link"]          =    "External link"; // value from english
//	$ARnls["ariadne:editor:hyperlinkedit"]          =    "Edit hyperlink"; // value from english
//	$ARnls["ariadne:editor:image_alttext"]          =    "Alternative text"; // value from english
//	$ARnls["ariadne:editor:image_settings"]         =    "Image settings"; // value from english
//	$ARnls["ariadne:editor:imageedit"]              =    "Edit image"; // value from english
//	$ARnls["ariadne:editor:internal_link"]          =    "Internal link"; // value from english
//	$ARnls["ariadne:editor:language"]               =    "Language"; // value from english
//	$ARnls["ariadne:editor:newwindow"]              =    "Open in new window"; // value from english
//	$ARnls["ariadne:editor:popup"]                  =    "Open in popup"; // value from english
//	$ARnls["ariadne:editor:preview"]                =    "Preview"; // value from english
//	$ARnls["ariadne:editor:style"]                  =    "Style"; // value from english
//	$ARnls["ariadne:err:rewrite.no_input"]          =    "Geef eerst herschrijfinstructies op."; // value from english
	$ARnls["ariadne:explore"]                       =    "Utforska";
	$ARnls["ariadne:export"]                        =    "Exportera";
//	$ARnls["ariadne:file_uploaded"]                 =    "File"; // value from english
	$ARnls["ariadne:folders"]                       =    "Mappar";
//	$ARnls["ariadne:generate"]                      =    "Generate"; // value from english
//	$ARnls["ariadne:grantkey"]                      =    "Grant key"; // value from english
	$ARnls["ariadne:grants"]                        =    "S&auml;tt r&auml;ttigheter f&ouml;r ";
//	$ARnls["ariadne:grants:grants_explained"]       =    "Grants explained for "; // value from english
//	$ARnls["ariadne:grants:objects_with_grants"]    =    "Objects with grants configured"; // value from english
//	$ARnls["ariadne:grants:other_grants"]           =    "Other grants for "; // value from english
//	$ARnls["ariadne:grants:users_with_grants"]      =    "Users/groups with grants on: "; // value from english
	$ARnls["ariadne:help"]                          =    "Hj&auml;lp";
	$ARnls["ariadne:iconview"]                      =    "V&auml;lj Ikon-vy";
//	$ARnls["ariadne:id"]                            =    "ID"; // value from english
	$ARnls["ariadne:import"]                        =    "Importera";
	$ARnls["ariadne:info"]                          =    "Information";
	$ARnls["ariadne:language"]                      =    "S&auml;tt spr&aring;k f&ouml;r ";
	$ARnls["ariadne:large"]                         =    "Ikoner";
//	$ARnls["ariadne:lastmodified"]                  =    "Last modified"; // value from english
	$ARnls["ariadne:link"]                          =    "L&auml;nk ";
//	$ARnls["ariadne:lock:toggle_all"]               =    "Toggle all"; // value from english
//	$ARnls["ariadne:logoff"]                        =    "Log off"; // value from english
//	$ARnls["ariadne:mimetype"]                      =    "MIME Type"; // value from english
//	$ARnls["ariadne:mogrify"]                       =    "Mogrify"; // value from english
	$ARnls["ariadne:new"]                           =    "L&auml;gg till nytt objekt";
//	$ARnls["ariadne:new:add_language"]              =    "Add language"; // value from english
//	$ARnls["ariadne:new:autonumber"]                =    "Number automatically"; // value from english
//	$ARnls["ariadne:new:below"]                     =    "Directly below the current object"; // value from english
//	$ARnls["ariadne:new:beside"]                    =    "Next to the current object at the same level"; // value from english
//	$ARnls["ariadne:new:change_type"]               =    "Change type"; // value from english
//	$ARnls["ariadne:new:create_object"]             =    "Create Object"; // value from english
//	$ARnls["ariadne:new:default_language_data"]     =    "Data for the default language"; // value from english
//	$ARnls["ariadne:new:display_name"]              =    "Display name"; // value from english
//	$ARnls["ariadne:new:extralanguages"]            =    "Add data for other languages"; // value from english
//	$ARnls["ariadne:new:filename"]                  =    "Filename"; // value from english
//	$ARnls["ariadne:new:lettersnumbers"]            =    "Use letters and numbers, no spaces"; // value from english
//	$ARnls["ariadne:new:location"]                  =    "Location"; // value from english
//	$ARnls["ariadne:new:select_type"]               =    "Choose the type of object to create:"; // value from english
//	$ARnls["ariadne:new:show_all_types"]            =    "Show all available types"; // value from english
//	$ARnls["ariadne:next"]                          =    "Next"; // value from english
//	$ARnls["ariadne:no_adding_found"]               =    "You can not add objects here."; // value from english
//	$ARnls["ariadne:no_objects_found"]              =    "No objects found."; // value from english
//	$ARnls["ariadne:object:copied_object"]          =    " (Copy)"; // value from english
//	$ARnls["ariadne:options"]                       =    "Options"; // value from english
//	$ARnls["ariadne:override_typetree"]             =    "Override typetree settings"; // value from english
//	$ARnls["ariadne:pdms:cmis_pass"]                =    "CMIS password"; // value from english
//	$ARnls["ariadne:pdms:cmis_root"]                =    "CMSI repository root"; // value from english
//	$ARnls["ariadne:pdms:cmis_url"]                 =    "CMIS URL"; // value from english
//	$ARnls["ariadne:pdms:cmis_user"]                =    "CMIS username"; // value from english
//	$ARnls["ariadne:pdms:ftp_host"]                 =    "FTP host"; // value from english
//	$ARnls["ariadne:pdms:ftp_pass"]                 =    "FTP password"; // value from english
//	$ARnls["ariadne:pdms:ftp_port"]                 =    "FTP port (default 21)"; // value from english
//	$ARnls["ariadne:pdms:ftp_root"]                 =    "FTP repository root"; // value from english
//	$ARnls["ariadne:pdms:ftp_user"]                 =    "FTP username"; // value from english
//	$ARnls["ariadne:pdms:pdms_type"]                =    "DMS type"; // value from english
	$ARnls["ariadne:preferences"]                   =    "Egenskaper";
//	$ARnls["ariadne:prev"]                          =    "Previous"; // value from english
	$ARnls["ariadne:priority"]                      =    "S&auml;tt prioritet f&ouml;r ";
	$ARnls["ariadne:programmers_reference"]         =    "Programmers Reference";
//	$ARnls["ariadne:query"]                         =    "Query"; // value from english
//	$ARnls["ariadne:remove_file"]                   =    "Remove current file"; // value from english
	$ARnls["ariadne:rename"]                        =    "Byt namn ";
//	$ARnls["ariadne:rewrite"]                       =    "Rewrite content"; // value from english
//	$ARnls["ariadne:rewrite.newreference"]          =    "New path"; // value from english
//	$ARnls["ariadne:rewrite.newurl"]                =    "New URL"; // value from english
//	$ARnls["ariadne:rewrite.oldreference"]          =    "Old path"; // value from english
//	$ARnls["ariadne:rewrite.oldurl"]                =    "Old URL"; // value from english
//	$ARnls["ariadne:rewrite.references"]            =    "Rewrite path references"; // value from english
//	$ARnls["ariadne:rewrite.urls"]                  =    "Rewrite URLs"; // value from english
//	$ARnls["ariadne:rewriting"]                     =    "Rewriting"; // value from english
	$ARnls["ariadne:search"]                        =    "S&ouml;k";
//	$ARnls["ariadne:selectlanguage"]                =    "Select a different language"; // value from english
	$ARnls["ariadne:settings"]                      =    "Inst&auml;llningar";
	$ARnls["ariadne:shortcut"]                      =    "&auml;ndra genv&auml;g";
	$ARnls["ariadne:small"]                         =    "Lista";
//	$ARnls["ariadne:su"]                            =    "Switch user"; // value from english
//	$ARnls["ariadne:svn"]                           =    "SVN"; // value from english
//	$ARnls["ariadne:svn:added"]                     =    "Added"; // value from english
//	$ARnls["ariadne:svn:checkout"]                  =    "Checkout"; // value from english
//	$ARnls["ariadne:svn:checkout_recursive"]        =    "SVN Recursive Checkout"; // value from english
//	$ARnls["ariadne:svn:checkunder"]                =    "Checkunder"; // value from english
//	$ARnls["ariadne:svn:checkunder_recursive"]      =    "SVN Recursive Checkunder"; // value from english
//	$ARnls["ariadne:svn:commit"]                    =    "Commit"; // value from english
//	$ARnls["ariadne:svn:commit_recursive"]          =    "SVN Recursive Commit"; // value from english
//	$ARnls["ariadne:svn:config"]                    =    "Configure"; // value from english
//	$ARnls["ariadne:svn:conflict"]                  =    "Conflict"; // value from english
//	$ARnls["ariadne:svn:delete"]                    =    "Delete"; // value from english
//	$ARnls["ariadne:svn:deleteconfirm"]             =    "Are you sure you want to delete this template from SVN?"; // value from english
//	$ARnls["ariadne:svn:deleted"]                   =    "Deleted"; // value from english
//	$ARnls["ariadne:svn:diff"]                      =    "Diff"; // value from english
//	$ARnls["ariadne:svn:import"]                    =    "Import"; // value from english
//	$ARnls["ariadne:svn:import_recursive"]          =    "SVN Recursive Import"; // value from english
//	$ARnls["ariadne:svn:info"]                      =    "SVN Info"; // value from english
//	$ARnls["ariadne:svn:insubversion"]              =    "In subversion"; // value from english
//	$ARnls["ariadne:svn:message"]                   =    "Message"; // value from english
//	$ARnls["ariadne:svn:modified"]                  =    "Modified"; // value from english
//	$ARnls["ariadne:svn:nomod"]                     =    "No modifications"; // value from english
//	$ARnls["ariadne:svn:notworkingcopy"]            =    "Not a working copy"; // value from english
//	$ARnls["ariadne:svn:password"]                  =    "SVN password"; // value from english
//	$ARnls["ariadne:svn:repository"]                =    "SVN repository"; // value from english
//	$ARnls["ariadne:svn:repository_information"]    =    "Repository information"; // value from english
//	$ARnls["ariadne:svn:resolved"]                  =    "Resolved"; // value from english
//	$ARnls["ariadne:svn:revert"]                    =    "Revert"; // value from english
//	$ARnls["ariadne:svn:revision"]                  =    "SVN Revision"; // value from english
//	$ARnls["ariadne:svn:settings"]                  =    "SVN Settings"; // value from english
//	$ARnls["ariadne:svn:unsvn"]                     =    "Remove version control"; // value from english
//	$ARnls["ariadne:svn:update"]                    =    "Update"; // value from english
//	$ARnls["ariadne:svn:update_recursive"]          =    "SVN Recursive Update"; // value from english
//	$ARnls["ariadne:svn:username"]                  =    "SVN username"; // value from english
//	$ARnls["ariadne:template:char"]                 =    "Char"; // value from english
//	$ARnls["ariadne:template:col"]                  =    "Col"; // value from english
//	$ARnls["ariadne:template:private"]              =    "Private"; // value from english
//	$ARnls["ariadne:template:row"]                  =    "Row"; // value from english
//	$ARnls["ariadne:template_editor"]               =    "Template editor"; // value from english
//	$ARnls["ariadne:templateeditor:ace"]            =    "ACE"; // value from english
//	$ARnls["ariadne:templateeditor:textarea"]       =    "Textarea"; // value from english
	$ARnls["ariadne:templates"]                     =    "S&auml;tt mallar f&ouml;r ";
//	$ARnls["ariadne:too_many_objects_found"]        =    "Too many objects found."; // value from english
	$ARnls["ariadne:tutorials"]                     =    "V&auml;gledning";
//	$ARnls["ariadne:type"]                          =    "Type"; // value from english
	$ARnls["ariadne:types"]                         =    "S&auml;tt typtr&auml;d f&ouml;r ";
//	$ARnls["ariadne:types:paddressbook"]            =    "Addressbook"; // value from english
//	$ARnls["ariadne:types:particle"]                =    "Article"; // value from english
//	$ARnls["ariadne:types:pbookmark"]               =    "Bookmark"; // value from english
//	$ARnls["ariadne:types:pcalendar"]               =    "Calendar"; // value from english
//	$ARnls["ariadne:types:pcalitem"]                =    "Calendar Item"; // value from english
//	$ARnls["ariadne:types:pdir"]                    =    "Directory"; // value from english
//	$ARnls["ariadne:types:pdir.projects"]           =    "Projects Folder"; // value from english
//	$ARnls["ariadne:types:pdms"]                    =    "DMS connection"; // value from english
//	$ARnls["ariadne:types:pfile"]                   =    "File"; // value from english
//	$ARnls["ariadne:types:pgroup"]                  =    "Group"; // value from english
//	$ARnls["ariadne:types:pldapconnection"]         =    "LDAP Connection"; // value from english
//	$ARnls["ariadne:types:pnewspaper"]              =    "Newspaper"; // value from english
//	$ARnls["ariadne:types:pobject"]                 =    "Object"; // value from english
//	$ARnls["ariadne:types:porganization"]           =    "Organization"; // value from english
//	$ARnls["ariadne:types:ppage"]                   =    "Page"; // value from english
//	$ARnls["ariadne:types:pperson"]                 =    "Person"; // value from english
//	$ARnls["ariadne:types:pphoto"]                  =    "Photo"; // value from english
//	$ARnls["ariadne:types:pphotobook"]              =    "Photobook"; // value from english
//	$ARnls["ariadne:types:pprofile"]                =    "Profile"; // value from english
//	$ARnls["ariadne:types:pproject"]                =    "Project"; // value from english
//	$ARnls["ariadne:types:pscenario"]               =    "Scenario"; // value from english
//	$ARnls["ariadne:types:psearch"]                 =    "Search"; // value from english
//	$ARnls["ariadne:types:psection"]                =    "Section"; // value from english
//	$ARnls["ariadne:types:pshortcut"]               =    "Shortcut"; // value from english
//	$ARnls["ariadne:types:psite"]                   =    "Site"; // value from english
//	$ARnls["ariadne:types:puser"]                   =    "User"; // value from english
	$ARnls["ariadne:up"]                            =    "Upp";
//	$ARnls["ariadne:uploading"]                     =    "Uploading..."; // value from english
	$ARnls["ariadne:view"]                          =    "Visa";
	$ARnls["ariadne:viewweb"]                       =    "Visa webbsida ";
//	$ARnls["ariadne:vtype"]                         =    "Virtual"; // value from english
//	$ARnls["ariadne:workspace:commit_selected"]     =    "Commit selected"; // value from english
//	$ARnls["ariadne:workspace:create"]              =    "Created"; // value from english
//	$ARnls["ariadne:workspace:delete"]              =    "Deleted"; // value from english
//	$ARnls["ariadne:workspace:diff_selected"]       =    "Diff selected"; // value from english
//	$ARnls["ariadne:workspace:manage_workspace"]    =    "Manage workspace"; // value from english
//	$ARnls["ariadne:workspace:move"]                =    "Moved"; // value from english
//	$ARnls["ariadne:workspace:revert_selected"]     =    "Revert selected"; // value from english
//	$ARnls["ariadne:workspace:status"]              =    "Status"; // value from english
//	$ARnls["ariadne:workspace:update"]              =    "Updated"; // value from english
//	$ARnls["ariadne:workspace:workspace"]           =    "Workspace"; // value from english
	$ARnls["ariadne:wysiwyg_editor"]                =    "WYSIWYG editor";
//	$ARnls["err:customdatanameinuse"]               =    "this name is already in use."; // value from english
//	$ARnls["err:defaultlanguagenotavailable"]       =    "The chosen default language was not selected as an available language."; // value from english
//	$ARnls["err:no_add_on_target"]                  =    "Sorry, no &quot;add&quot; grants on target"; // value from english
//	$ARnls["err:nocustomdataname"]                  =    "You must enter a name."; // value from english
//	$ARnls["err:nosalt"]                            =    "No salt is configured in Ariadne. Please configure this in the main Ariadne configuration to allow generation of grant keys."; // value from english
//	$ARnls["err:svn:enterURL"]                      =    "Please enter a valid SVN repository URL."; // value from english
//	$ARnls["err:svn:leaving_recurse_tree"]          =    "This repository is not part of the repository tree of the parent."; // value from english
//	$ARnls["err:typetree_does_not_allow"]           =    "Typetree does not allow this object type here"; // value from english


?>