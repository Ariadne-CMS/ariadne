<?php


	/*****************************************************************************

		The Swedish nls files are contributed by: Niklas Koskela <ntkk@htc.se>
                                                      Karl Thysell <karl@htc.se>

	*****************************************************************************/

	$ARnls["ariadne:about"]						=	"Om...";
	$ARnls["ariadne:browsebydate"]				=	"Bl&auml;ddra per datum";
	$ARnls["ariadne:browsebyletter"]				=	"Bl&auml;ddra per bokstav";
	$ARnls["ariadne:cache"]						=	"S&auml;tt cache f&ouml;r ";
	$ARnls["ariadne:copy"]						=	"Kopiera ";
	$ARnls["ariadne:customfields"]				=	"S&auml;tt anpassade f&auml;lt f&ouml;r ";
	$ARnls["ariadne:delete"]						=	"Radera ";
	$ARnls["ariadne:details"]					=	"Detaljer";
	$ARnls["ariadne:detailsH"]					=	"Mera...";
	$ARnls["ariadne:edit"]						=	"&auml;ndra ";
	$ARnls["ariadne:explore"]					=	"Utforska";
	$ARnls["ariadne:export"]						=	"Exportera";
	$ARnls["ariadne:folders"]					=	"Mappar";
	$ARnls["ariadne:grants"]						=	"S&auml;tt r&auml;ttigheter f&ouml;r ";
	$ARnls["ariadne:help"]						=	"Hj&auml;lp";
	$ARnls["ariadne:iconview"]					=	"V&auml;lj Ikon-vy";
	$ARnls["ariadne:import"]						=	"Importera";
	$ARnls["ariadne:info"]						=	"Information";
	$ARnls["ariadne:language"]					=	"S&auml;tt spr&aring;k f&ouml;r ";
	$ARnls["ariadne:large"]						=	"Ikoner";
	$ARnls["ariadne:link"]						=	"L&auml;nk ";
	$ARnls["ariadne:new"]						=	"L&auml;gg till nytt objekt";
	$ARnls["ariadne:preferences"]				=	"Egenskaper";
	$ARnls["ariadne:priority"]					=	"S&auml;tt prioritet f&ouml;r ";
	$ARnls["ariadne:rename"]						=	"Byt namn ";
	$ARnls["ariadne:search"]						=	"S&ouml;k";
	$ARnls["ariadne:settings"]					=	"Inst&auml;llningar";
	$ARnls["ariadne:shortcut"]					=	"&auml;ndra genv&auml;g";
	$ARnls["ariadne:small"]						=	"Lista";
	$ARnls["ariadne:templates"]					=	"S&auml;tt mallar f&ouml;r ";
	$ARnls["ariadne:tutorials"]					=	"V&auml;gledning";
	$ARnls["ariadne:types"]						=	"S&auml;tt typtr&auml;d f&ouml;r ";
	$ARnls["ariadne:up"]							=	"Upp";
	$ARnls["ariadne:view"]						=	"Visa";
	$ARnls["ariadne:viewweb"]					=	"Visa webbsida ";
	$ARnls['ariadne:wysiwyg_editor']			=	"WYSIWYG editor";

	$ARnls['ariadne:programmers_reference']		= 'Programmers Reference';
	$ARnls['ariadne:ace_editor']				= 'Ace Editor';

?>